Photodiode Amplifier Circuit


.include ua741.txt
.include Diode_1N914.txt
.include zener_1N4732A.txt


x1 1 2 3 4 5 UA741
r2 3 7 13.3k
r1 4 8 13.3k
vcc 3 0 15
vdd 4 0 -15
vin 2 0 
d1 7 5 1N914
d2 7 6 1N914
d3 5 8 1N914
d4 6 8 1N914
x2 6 9 DI_1N4732A
x3 0 9 DI_1N4732A
vdummy 1 6 0

.dc vin 10 -10 0.1

.control

run

plot v(1)

.endc
.end