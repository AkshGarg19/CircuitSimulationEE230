Photodiode Amplifier Circuit


.include lm324.txt


x1 1 2 3 4 5 LM324
r2 6 8 10.1k
r1 8 0 9.5k
rg 2 7 9.8k
rf 2 5 164.8k
vcc 3 0 5
vdd 4 0 0
vin 7 0 
vref 6 0 1.22
vos 1 8 2m

.dc vin 0 2 2m

.control

run

plot v(5)

.endc
.end